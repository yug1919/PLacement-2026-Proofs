library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity FDE is
port(clk, reset: in std_logic;
	  opcode : in std_logic_vector(3 downto 0);
     lsb : in std_logic_vector(2 downto 0);
	  cont_signal : out std_logic_vector(31 downto 0));
end entity FDE;

architecture contr of FDE is
    signal C0_2, C0_3, C1_4, C0_4, C1_5, C0_5, C0_11, C0_6, C1_6, C2_7, C1_7, C0_7,
	 C1_A1, C0_A1, C1_W, Z1_W, C1_8, C0_8, C1_9, C0_9, C1_A3,
	 C0_A3, C_W, Z_W, C0_10, DMEM_W, DMEM_M, IS_NONE, IS_CEC1,
	 IP_W, RF_W, RF_M: std_logic;

	 
begin

reset_proc: process(reset)
begin
if (reset = '1') then
	C0_2    <= '0';
	C0_3    <= '0';
	C1_4    <= '0';
	C0_4    <= '0';
	C1_5    <= '0';
	C0_5    <= '0';
	C0_11   <= '0';
	C1_6    <= '0';
	C0_6    <= '0';
	C2_7    <= '0';
	C1_7    <= '0';
	C0_7    <= '0';
	C1_A1   <= '0';
	C0_A1   <= '0';
	C1_W    <= '0';
	Z1_W    <= '0';
	C1_8    <= '0';
	C0_8    <= '0';
	C1_9    <= '0';
	C0_9    <= '0';
	C1_A3   <= '0';
	C0_A3   <= '0';
	C_W     <= '0';
	Z_W     <= '0';
	C0_10   <= '0';
	DMEM_W  <= '0';
	DMEM_M  <= '0';
	IS_NONE <= '0';
	IS_CEC1 <= '0';
	IP_W    <= '0';
	RF_W    <= '0';
	RF_M    <= '0';
end if;
end process reset_proc;
    control_check: process(opcode, lsb, clk)
    begin
        
        C0_2 <= '0';
        C0_3 <= '0';
        C1_4 <= '0';
        C0_4 <= '0';
        C1_5 <= '0';
        C0_5 <= '0';
		  C0_11 <= '0';
        C1_6 <= '0';
        C0_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '0';
        C0_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '0';
        C0_8 <= '0';
        C1_9 <= '0';
        C0_9 <= '0';
        C1_A3 <= '0';
        C0_A3 <= '0';
        C_W <= '0';
        Z_W <= '0';
        C0_10 <= '0';
        DMEM_W <= '0';
        DMEM_M <= '0';
        IS_NONE <= '0';
        IS_CEC1 <= '0';
        IP_W <= '0';
        RF_W <= '0';
        RF_M <= '0';
     
        case opcode is
            when "0000" =>
                C0_2 <= '1';
                C0_3 <= '0';
                C1_4 <= '0';
                C0_4 <= '1';
                C1_5 <= '1';
                C0_5 <= '0';
                C0_6 <= '0';
					 C1_6 <= '0';
                C2_7 <= '0';
                C1_7 <= '1';
                C0_7 <= '0';
                C1_A1 <= '0';
                C0_A1 <= '0';
                C1_W <= '1';
                Z1_W <= '1';
                C1_8 <= '1';
                C0_8 <= '0';
                C1_9 <= '1';
                C0_9 <= '1';
                C1_A3 <= '1';
                C0_A3 <= '1';
                C_W <= '1';
                Z_W <= '1';
                IS_NONE <= '1';
                IS_CEC1 <= '1';
                IP_W <= '1';
                RF_W <= '1';
                RF_M <= '0';
            when "0001" =>
				case lsb is
				when "000" | "010" | "001" | "100" | "110" | "101" =>
        C0_2 <= '1';
        C0_3 <= '1';
        C1_4 <= '0';
        C0_4 <= '0';
        C1_5 <= '1';
        C0_5 <= '0';
        C0_6 <= '0';
        C1_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '1';
        Z1_W <= '1';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '1';
        Z_W <= '1';
        IS_NONE <= '1';
        IS_CEC1 <= '1';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
		   if (lsb = "000") or (lsb = "010") or (lsb = "001") then
			  C0_7 <= '0';
			  
			elsif (lsb = "100") or (lsb = "110") or (lsb = "101") then
			  C0_7 <= '1';
			  
			 end if;
			 
			when "011" | "111" =>
		  C0_2 <= '1';
        C0_3 <= '1';
        C1_4 <= '0';
        C0_4 <= '0';
        C1_5 <= '0';
        C0_5 <= '0';
		  C0_11 <= '1';
        C0_6 <= '0';
        C1_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '0';
        C0_8 <= '0';
        C1_9 <= '0';
        C0_9 <= '0';
        C1_A3 <= '0';
        C0_A3 <= '0';
        C_W <= '1';
        Z_W <= '1';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
			if (lsb = "011") then
			  C0_7 <= '0';
			  
			elsif (lsb = "111") then
			  C0_7 <= '1';
			  
			 end if; 
			 
			 end case;
			 
			when "0010" =>
		  C0_2 <= '1';
        C0_3 <= '1';
        C1_4 <= '0';
        C0_4 <= '0';
        C1_5 <= '1';
        C0_5 <= '0';
        C0_6 <= '0';
        C1_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '1';
        C1_W <= '1';
        Z1_W <= '1';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '1';
        Z_W <= '1';
        IS_NONE <= '1';
        IS_CEC1 <= '1';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
			 
			  if (lsb = "000") or (lsb = "010") or (lsb = "001") then
			  C0_7 <= '0';
			  
			elsif (lsb = "100") or (lsb = "110") or (lsb = "101") then
			  C0_7 <= '1';
			  
			  end if;
			  
         
            when "0011" =>
        C0_2 <= '0';
        C0_3 <= '0';
        C1_4 <= '1';
        C0_4 <= '0';
        C1_5 <= '0';
        C0_5 <= '0';
		  C0_11 <= '0';
        C1_6 <= '0';
        C0_6 <= '1';
        C2_7 <= '1';
        C1_7 <= '0';
		  C0_7 <= '0';
        C1_A1 <= '1';
        C0_A1 <= '1';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
		  
		  when "0100" =>
        C0_2 <= '0';
        C0_3 <= '1';
        C1_4 <= '1';
        C0_4 <= '0';
        C1_5 <= '1';
        C0_5 <= '0';
        C1_6 <= '1';
        C0_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '1';
		  C0_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '1';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '1';
		  C0_10 <= '0';
		  DMEM_W <= '0';
		  DMEM_M <= '0';
        IS_NONE <= '0';
        IS_CEC1 <= '1';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
		  
		  when "0101" =>
        C0_2 <= '1';
        C0_3 <= '1';
        C1_6 <= '1';
        C0_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '1';
		  C0_7 <= '0';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
		  C0_10 <= '0';
		  DMEM_W <= '1';
		  DMEM_M <= '0';
        IS_NONE <= '0';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '0';
        RF_M <= '0';
		  
		   when "0110" =>
        C0_2 <= '1';
        C0_3 <= '0';
        C1_6 <= '0';
        C0_6 <= '1';
        C2_7 <= '1';
        C1_7 <= '0';
        C0_7 <= '0';
        C1_A1 <= '1';
        C0_A1 <= '1';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
        C0_10 <= '1';
        DMEM_W <= '0';
        DMEM_M <= '1';
        IS_NONE <= '0';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '1';
		  
		  when "0111" =>
        C0_2 <= '1';
        C0_3 <= '0';
        C1_6 <= '0';
        C0_6 <= '1';
        C2_7 <= '1';
        C1_7 <= '0';
        C0_7 <= '0';
        C1_A1 <= '1';
        C0_A1 <= '1';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
        C0_10 <= '1';
        DMEM_W <= '1';
        DMEM_M <= '1';
        IS_NONE <= '0';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '0';
        RF_M <= '1';
     
	     when "1000" | "1001" =>
	     C0_2 <= '1';
        C0_3 <= '1';
        C1_6 <= '0';
        C0_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '0';
        C0_7 <= '0';
        C1_A1 <= '1';
        C0_A1 <= '0';
        C1_W <= '1';
        Z1_W <= '1';
        C1_8 <= '0';
        C0_8 <= '1';
        C1_9 <= '0';
        C0_9 <= '1';
        C1_A3 <= '0';
        C0_A3 <= '0';
        C_W <= '0';
        Z_W <= '0';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '0';
        RF_M <= '0';
		  
		  when "1100" =>
		  C0_2 <= '0';
        C0_3 <= '0';
        C1_4 <= '1';
        C0_4 <= '0';
        C1_5 <= '1';
        C0_5 <= '0';
		  C0_11 <= '1';
        C1_6 <= '1';
        C0_6 <= '1';
        C2_7 <= '1';
        C1_7 <= '0';
        C0_7 <= '1';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '0';
        C0_8 <= '1';
        C1_9 <= '1';
        C0_9 <= '0';
        C1_A3 <= '0';
        C0_A3 <= '0';
        C_W <= '0';
        Z_W <= '0';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
		 
		  when "1101" =>
		  
		  C0_2 <= '0';
        C0_3 <= '1';
        C1_4 <= '1';
        C0_4 <= '0';
        C1_5 <= '1';
        C0_5 <= '0';
        C1_6 <= '1';
        C0_6 <= '1';
        C2_7 <= '1';
        C1_7 <= '0';
        C0_7 <= '1';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '1';
        RF_M <= '0';
		   
		when "1111" =>
		  C0_2 <= '1';
        C0_3 <= '0';
        C1_6 <= '0';
        C0_6 <= '0';
        C2_7 <= '0';
        C1_7 <= '1';
        C0_7 <= '1';
        C1_A1 <= '0';
        C0_A1 <= '0';
        C1_W <= '0';
        Z1_W <= '0';
        C1_8 <= '1';
        C0_8 <= '0';
        C1_9 <= '1';
        C0_9 <= '1';
        C1_A3 <= '1';
        C0_A3 <= '1';
        C_W <= '0';
        Z_W <= '0';
        IS_NONE <= '1';
        IS_CEC1 <= '0';
        IP_W <= '1';
        RF_W <= '0';
        RF_M <= '0';
               
            when others =>
                null;
        end case;

    end process;
end contr;
